package keccak_testbench_pkg;
  import uvm_pkg::*;
  
  `include "keccak_sequence.sv"
  `include "keccak_driver.sv"
  `include "keccak_monitor.sv"
  `include "keccak_scoreboard.sv"

  //Include subscriber to package
    `include "keccak_subscriber.sv"

  `include "keccak_agent.sv"
  `include "keccak_env.sv"
  `include "keccak_test.sv"

endpackage
  
